library verilog;
use verilog.vl_types.all;
entity tbCompressor is
end tbCompressor;
