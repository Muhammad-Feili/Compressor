library verilog;
use verilog.vl_types.all;
entity tbComp5to1 is
end tbComp5to1;
